module Mul3 (in_byte,out_byte);
    input [7:0] in_byte;
    output reg [7:0] out_byte;

    reg [7:0] Mul3_Table [0:255];
    
initial begin
    Mul3_Table[0]   = 8'h00;
    Mul3_Table[1]   = 8'h03;
    Mul3_Table[2]   = 8'h06;
    Mul3_Table[3]   = 8'h05;
    Mul3_Table[4]   = 8'h0c;
    Mul3_Table[5]   = 8'h0f;
    Mul3_Table[6]   = 8'h0a;
    Mul3_Table[7]   = 8'h09;
    Mul3_Table[8]   = 8'h18;
    Mul3_Table[9]   = 8'h1b;
    Mul3_Table[10]  = 8'h1e;
    Mul3_Table[11]  = 8'h1d;
    Mul3_Table[12]  = 8'h14;
    Mul3_Table[13]  = 8'h17;
    Mul3_Table[14]  = 8'h12;
    Mul3_Table[15]  = 8'h11;
    Mul3_Table[16]  = 8'h30;
    Mul3_Table[17]  = 8'h33;
    Mul3_Table[18]  = 8'h36;
    Mul3_Table[19]  = 8'h35;
    Mul3_Table[20]  = 8'h3c;
    Mul3_Table[21]  = 8'h3f;
    Mul3_Table[22]  = 8'h3a;
    Mul3_Table[23]  = 8'h39;
    Mul3_Table[24]  = 8'h28;
    Mul3_Table[25]  = 8'h2b;
    Mul3_Table[26]  = 8'h2e;
    Mul3_Table[27]  = 8'h2d;
    Mul3_Table[28]  = 8'h24;
    Mul3_Table[29]  = 8'h27;
    Mul3_Table[30]  = 8'h22;
    Mul3_Table[31]  = 8'h21;
    Mul3_Table[32]  = 8'h60;
    Mul3_Table[33]  = 8'h63;
    Mul3_Table[34]  = 8'h66;
    Mul3_Table[35]  = 8'h65;
    Mul3_Table[36]  = 8'h6c;
    Mul3_Table[37]  = 8'h6f;
    Mul3_Table[38]  = 8'h6a;
    Mul3_Table[39]  = 8'h69;
    Mul3_Table[40]  = 8'h78;
    Mul3_Table[41]  = 8'h7b;
    Mul3_Table[42]  = 8'h7e;
    Mul3_Table[43]  = 8'h7d;
    Mul3_Table[44]  = 8'h74;
    Mul3_Table[45]  = 8'h77;
    Mul3_Table[46]  = 8'h72;
    Mul3_Table[47]  = 8'h71;
    Mul3_Table[48]  = 8'h50;
    Mul3_Table[49]  = 8'h53;
    Mul3_Table[50]  = 8'h56;
    Mul3_Table[51]  = 8'h55;
    Mul3_Table[52]  = 8'h5c;
    Mul3_Table[53]  = 8'h5f;
    Mul3_Table[54]  = 8'h5a;
    Mul3_Table[55]  = 8'h59;
    Mul3_Table[56]  = 8'h48;
    Mul3_Table[57]  = 8'h4b;
    Mul3_Table[58]  = 8'h4e;
    Mul3_Table[59]  = 8'h4d;
    Mul3_Table[60]  = 8'h44;
    Mul3_Table[61]  = 8'h47;
    Mul3_Table[62]  = 8'h42;
    Mul3_Table[63]  = 8'h41;
    Mul3_Table[64]  = 8'hc0;
    Mul3_Table[65]  = 8'hc3;
    Mul3_Table[66]  = 8'hc6;
    Mul3_Table[67]  = 8'hc5;
    Mul3_Table[68]  = 8'hcc;
    Mul3_Table[69]  = 8'hcf;
    Mul3_Table[70]  = 8'hca;
    Mul3_Table[71]  = 8'hc9;
    Mul3_Table[72]  = 8'hd8;
    Mul3_Table[73]  = 8'hdb;
    Mul3_Table[74]  = 8'hde;
    Mul3_Table[75]  = 8'hdd;
    Mul3_Table[76]  = 8'hd4;
    Mul3_Table[77]  = 8'hd7;
    Mul3_Table[78]  = 8'hd2;
Mul3_Table[79]  = 8'hd1;
Mul3_Table[80]  = 8'hf0;
Mul3_Table[81]  = 8'hf3;
Mul3_Table[82]  = 8'hf6;
Mul3_Table[83]  = 8'hf5;
Mul3_Table[84]  = 8'hfc;
Mul3_Table[85]  = 8'hff;
Mul3_Table[86]  = 8'hfa;
Mul3_Table[87]  = 8'hf9;
Mul3_Table[88]  = 8'he8;
Mul3_Table[89]  = 8'heb;
Mul3_Table[90]  = 8'hee;
Mul3_Table[91]  = 8'hed;
Mul3_Table[92]  = 8'he4;
Mul3_Table[93]  = 8'he7;
Mul3_Table[94]  = 8'he2;
Mul3_Table[95]  = 8'he1;
Mul3_Table[96]  = 8'ha0;
Mul3_Table[97]  = 8'ha3;
Mul3_Table[98]  = 8'ha6;
Mul3_Table[99]  = 8'ha5;
Mul3_Table[100] = 8'hac;
Mul3_Table[101] = 8'haf;
Mul3_Table[102] = 8'haa;
Mul3_Table[103] = 8'ha9;
Mul3_Table[104] = 8'hb8;
Mul3_Table[105] = 8'hbb;
Mul3_Table[106] = 8'hbe;
Mul3_Table[107] = 8'hbd;
Mul3_Table[108] = 8'hb4;
Mul3_Table[109] = 8'hb7;
Mul3_Table[110] = 8'hb2;
Mul3_Table[111] = 8'hb1;
Mul3_Table[112] = 8'h90;
Mul3_Table[113] = 8'h93;
Mul3_Table[114] = 8'h96;
Mul3_Table[115] = 8'h95;
Mul3_Table[116] = 8'h9c;
Mul3_Table[117] = 8'h9f;
Mul3_Table[118] = 8'h9a;
Mul3_Table[119] = 8'h99;
Mul3_Table[120] = 8'h88;
Mul3_Table[121] = 8'h8b;
Mul3_Table[122] = 8'h8e;
Mul3_Table[123] = 8'h8d;
Mul3_Table[124] = 8'h84;
Mul3_Table[125] = 8'h87;
Mul3_Table[126] = 8'h82;
Mul3_Table[127] = 8'h81;
Mul3_Table[128] = 8'h9b;
Mul3_Table[129] = 8'h98;
Mul3_Table[130] = 8'h9d;
Mul3_Table[131] = 8'h9e;
Mul3_Table[132] = 8'h97;
Mul3_Table[133] = 8'h94;
Mul3_Table[134] = 8'h91;
Mul3_Table[135] = 8'h92;
Mul3_Table[136] = 8'h83;
Mul3_Table[137] = 8'h80;
Mul3_Table[138] = 8'h85;
Mul3_Table[139] = 8'h86;
Mul3_Table[140] = 8'h8f;
Mul3_Table[141] = 8'h8c;
Mul3_Table[142] = 8'h89;
Mul3_Table[143] = 8'h8a;
Mul3_Table[144] = 8'hab;
Mul3_Table[145] = 8'ha8;
Mul3_Table[146] = 8'had;
  Mul3_Table[147] = 8'hae; Mul3_Table[148] = 8'ha7; Mul3_Table[149] = 8'ha4; Mul3_Table[150] = 8'ha1;
  Mul3_Table[151] = 8'ha2; Mul3_Table[152] = 8'hb3; Mul3_Table[153] = 8'hb0; Mul3_Table[154] = 8'hb5;
  Mul3_Table[155] = 8'hb6; Mul3_Table[156] = 8'hbf; Mul3_Table[157] = 8'hbc; Mul3_Table[158] = 8'hb9;
  Mul3_Table[159] = 8'hba; Mul3_Table[160] = 8'hfb; Mul3_Table[161] = 8'hf8; Mul3_Table[162] = 8'hfd;
  Mul3_Table[163] = 8'hfe; Mul3_Table[164] = 8'hf7; Mul3_Table[165] = 8'hf4; Mul3_Table[166] = 8'hf1;
  Mul3_Table[167] = 8'hf2; Mul3_Table[168] = 8'he3; Mul3_Table[169] = 8'he0; Mul3_Table[170] = 8'he5;
  Mul3_Table[171] = 8'he6; Mul3_Table[172] = 8'hef; Mul3_Table[173] = 8'hec; Mul3_Table[174] = 8'he9;
  Mul3_Table[175] = 8'hea; Mul3_Table[176] = 8'hcb; Mul3_Table[177] = 8'hc8; Mul3_Table[178] = 8'hcd;
  Mul3_Table[179] = 8'hce; Mul3_Table[180] = 8'hc7; Mul3_Table[181] = 8'hc4; Mul3_Table[182] = 8'hc1;
  Mul3_Table[183] = 8'hc2; Mul3_Table[184] = 8'hd3; Mul3_Table[185] = 8'hd0; Mul3_Table[186] = 8'hd5;
  Mul3_Table[187] = 8'hd6; Mul3_Table[188] = 8'hdf; Mul3_Table[189] = 8'hdc; Mul3_Table[190] = 8'hd9;
  Mul3_Table[191] = 8'hda; Mul3_Table[192] = 8'h5b; Mul3_Table[193] = 8'h58; Mul3_Table[194] = 8'h5d;
  Mul3_Table[195] = 8'h5e; Mul3_Table[196] = 8'h57; Mul3_Table[197] = 8'h54; Mul3_Table[198] = 8'h51;
  Mul3_Table[199] = 8'h52; Mul3_Table[200] = 8'h43; Mul3_Table[201] = 8'h40; Mul3_Table[202] = 8'h45;
  Mul3_Table[203] = 8'h46; Mul3_Table[204] = 8'h4f; Mul3_Table[205] = 8'h4c; Mul3_Table[206] = 8'h49;
  Mul3_Table[207] = 8'h4a; Mul3_Table[208] = 8'h6b; Mul3_Table[209] = 8'h68; Mul3_Table[210] = 8'h6d;
  Mul3_Table[211] = 8'h6e; Mul3_Table[212] = 8'h67; Mul3_Table[213] = 8'h64; Mul3_Table[214] = 8'h61;
  Mul3_Table[215] = 8'h62; Mul3_Table[216] = 8'h73; Mul3_Table[217] = 8'h70; Mul3_Table[218] = 8'h75;
  Mul3_Table[219] = 8'h76; Mul3_Table[220] = 8'h7f; Mul3_Table[221] = 8'h7c; Mul3_Table[222] = 8'h79;
  Mul3_Table[223] = 8'h7a; Mul3_Table[224] = 8'h3b; Mul3_Table[225] = 8'h38; Mul3_Table[226] = 8'h3d;
  Mul3_Table[227] = 8'h3e; Mul3_Table[228] = 8'h37; Mul3_Table[229] = 8'h34; Mul3_Table[230] = 8'h31;
  Mul3_Table[231] = 8'h32; Mul3_Table[232] = 8'h23; Mul3_Table[233] = 8'h20; Mul3_Table[234] = 8'h25;
  Mul3_Table[235] = 8'h26; Mul3_Table[236] = 8'h2f; Mul3_Table[237] = 8'h2c; Mul3_Table[238] = 8'h29;
  Mul3_Table[239] = 8'h2a; Mul3_Table[240] = 8'h0b; Mul3_Table[241] = 8'h08; Mul3_Table[242] = 8'h0d;
  Mul3_Table[243] = 8'h0e; Mul3_Table[244] = 8'h07; Mul3_Table[245] = 8'h04; Mul3_Table[246] = 8'h01;
  Mul3_Table[247] = 8'h02; Mul3_Table[248] = 8'h13; Mul3_Table[249] = 8'h10; Mul3_Table[250] = 8'h15;
  Mul3_Table[251] = 8'h16; Mul3_Table[252] = 8'h1f; Mul3_Table[253] = 8'h1c; Mul3_Table[254] = 8'h19;
  Mul3_Table[255] = 8'h1a;
end

    assign out_byte = Mul3_Table[in_byte];

endmodule